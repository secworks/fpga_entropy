
module inv1(
            input wire  s,
            output wire d
           );


  assign d = ~s;
  
endmodule // inv1

  
